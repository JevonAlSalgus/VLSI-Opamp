magic
tech sky130A
magscale 1 2
timestamp 1729268141
<< nwell >>
rect -243 -1747 582 535
<< nsubdiff >>
rect -207 465 -151 499
rect 490 465 546 499
rect -207 439 -173 465
rect 512 439 546 465
rect -207 -1677 -173 -1651
rect 512 -1677 546 -1651
rect -207 -1711 -151 -1677
rect 490 -1711 546 -1677
<< nsubdiffcont >>
rect -151 465 490 499
rect -207 -1651 -173 439
rect 512 -1651 546 439
rect -151 -1711 490 -1677
<< poly >>
rect -47 16 -17 47
rect -109 0 -17 16
rect -109 -34 -93 0
rect -59 -34 -17 0
rect -109 -50 -17 -34
rect 357 16 387 47
rect 357 0 449 16
rect 357 -34 399 0
rect 433 -34 449 0
rect 357 -50 449 -34
rect -47 -484 -17 -453
rect -109 -500 -17 -484
rect -109 -534 -93 -500
rect -59 -534 -17 -500
rect -109 -550 -17 -534
rect 357 -484 387 -453
rect 357 -500 449 -484
rect 357 -534 399 -500
rect 433 -534 449 -500
rect 357 -550 449 -534
rect -109 -672 -17 -656
rect 41 -657 141 -550
rect 199 -657 299 -550
rect -109 -706 -93 -672
rect -59 -706 -17 -672
rect -109 -722 -17 -706
rect -47 -753 -17 -722
rect 357 -672 449 -656
rect 357 -706 399 -672
rect 433 -706 449 -672
rect 357 -722 449 -706
rect 357 -753 387 -722
rect -109 -1172 -17 -1156
rect -109 -1206 -93 -1172
rect -59 -1206 -17 -1172
rect -109 -1222 -17 -1206
rect -47 -1253 -17 -1222
rect 357 -1172 449 -1156
rect 357 -1206 399 -1172
rect 433 -1206 449 -1172
rect 357 -1222 449 -1206
rect 357 -1253 387 -1222
<< polycont >>
rect -93 -34 -59 0
rect 399 -34 433 0
rect -93 -534 -59 -500
rect 399 -534 433 -500
rect -93 -706 -59 -672
rect 399 -706 433 -672
rect -93 -1206 -59 -1172
rect 399 -1206 433 -1172
<< locali >>
rect -207 465 -151 499
rect 490 465 546 499
rect -207 439 -173 465
rect 512 439 546 465
rect -93 0 -59 47
rect 399 0 433 59
rect -109 -34 -93 0
rect -59 -34 -43 0
rect 383 -34 399 0
rect 433 -34 449 0
rect -93 -500 -59 -453
rect 399 -500 433 -453
rect -109 -534 -93 -500
rect -59 -534 -43 -500
rect 383 -534 399 -500
rect 433 -534 449 -500
rect -109 -706 -93 -672
rect -59 -706 -43 -672
rect 383 -706 399 -672
rect 433 -706 449 -672
rect -93 -753 -59 -706
rect 399 -753 433 -706
rect -109 -1206 -93 -1172
rect -59 -1206 -43 -1172
rect 383 -1206 399 -1172
rect 433 -1206 449 -1172
rect -93 -1253 -59 -1206
rect 399 -1253 433 -1206
rect -207 -1677 -173 -1651
rect 512 -1677 546 -1651
rect -207 -1711 -151 -1677
rect 490 -1711 546 -1677
<< viali >>
rect 57 465 125 499
rect -93 -34 -59 0
rect 399 -34 433 0
rect -93 -534 -59 -500
rect 399 -534 433 -500
rect -93 -706 -59 -672
rect 399 -706 433 -672
rect -93 -1206 -59 -1172
rect 399 -1206 433 -1172
<< metal1 >>
rect 45 499 137 505
rect 45 465 57 499
rect 125 465 137 499
rect 45 459 137 465
rect -59 235 -5 247
rect -112 59 -102 235
rect -50 59 29 235
rect 134 59 144 235
rect 196 59 206 235
rect 292 59 302 235
rect 354 59 433 235
rect -99 6 -53 47
rect -105 0 -47 6
rect -105 -34 -93 0
rect -59 -34 -47 0
rect -105 -40 -47 -34
rect 57 -89 125 -34
rect 205 -43 215 9
rect 283 -43 293 9
rect 393 6 439 59
rect 387 0 445 6
rect 387 -34 399 0
rect 433 -34 445 0
rect 387 -40 445 -34
rect 57 -131 283 -89
rect 47 -215 57 -163
rect 125 -215 135 -163
rect 215 -172 283 -131
rect -93 -441 -14 -265
rect 38 -441 48 -265
rect 134 -441 144 -265
rect 196 -441 206 -265
rect 311 -441 390 -265
rect 442 -441 452 -265
rect -99 -494 -53 -453
rect 393 -494 439 -453
rect -105 -500 -47 -494
rect -105 -534 -93 -500
rect -59 -534 -47 -500
rect -105 -540 -47 -534
rect 387 -500 445 -494
rect 387 -534 399 -500
rect 433 -534 445 -500
rect 387 -540 445 -534
rect -105 -672 -47 -666
rect -105 -706 -93 -672
rect -59 -706 -47 -672
rect -105 -712 -47 -706
rect 387 -672 445 -666
rect 387 -706 399 -672
rect 433 -706 445 -672
rect 387 -712 445 -706
rect -99 -753 -53 -712
rect 393 -753 439 -712
rect -93 -941 -14 -765
rect 38 -941 48 -765
rect 134 -941 144 -765
rect 196 -941 206 -765
rect 311 -941 390 -765
rect 442 -941 452 -765
rect 47 -1043 57 -991
rect 125 -1043 135 -991
rect 215 -1081 283 -1034
rect 57 -1123 283 -1081
rect -105 -1172 -47 -1166
rect 57 -1172 125 -1123
rect -105 -1206 -93 -1172
rect -59 -1206 -47 -1172
rect -105 -1212 -47 -1206
rect -99 -1253 -53 -1212
rect 205 -1215 215 -1163
rect 283 -1215 293 -1163
rect 387 -1172 445 -1166
rect 387 -1206 399 -1172
rect 433 -1206 445 -1172
rect 387 -1212 445 -1206
rect 393 -1253 439 -1212
rect -112 -1441 -102 -1265
rect -50 -1441 29 -1265
rect 134 -1441 144 -1265
rect 196 -1441 206 -1265
rect 292 -1441 302 -1265
rect 354 -1441 433 -1265
<< via1 >>
rect -102 59 -50 235
rect 144 59 196 235
rect 302 59 354 235
rect 215 -43 283 9
rect 57 -215 125 -163
rect -14 -441 38 -265
rect 144 -441 196 -265
rect 390 -441 442 -265
rect -14 -941 38 -765
rect 144 -941 196 -765
rect 390 -941 442 -765
rect 57 -1043 125 -991
rect 215 -1215 283 -1163
rect -102 -1441 -50 -1265
rect 144 -1441 196 -1265
rect 302 -1441 354 -1265
<< metal2 >>
rect -5 347 345 376
rect -104 235 -48 245
rect -104 49 -48 59
rect -5 -255 29 347
rect 311 245 345 347
rect 142 235 198 245
rect 142 49 198 59
rect 302 235 354 245
rect 302 49 354 59
rect 215 9 283 19
rect 215 -89 283 -43
rect 57 -138 283 -89
rect 57 -163 125 -138
rect 57 -225 125 -215
rect -14 -265 38 -255
rect -14 -451 38 -441
rect 142 -265 198 -255
rect 142 -451 198 -441
rect -5 -755 29 -451
rect -14 -765 38 -755
rect -14 -951 38 -941
rect 142 -765 198 -755
rect 142 -951 198 -941
rect -104 -1265 -48 -1255
rect -104 -1451 -48 -1441
rect -5 -1553 29 -951
rect 57 -991 125 -981
rect 57 -1081 125 -1043
rect 57 -1130 283 -1081
rect 215 -1163 283 -1130
rect 215 -1225 283 -1215
rect 311 -1255 345 49
rect 388 -265 444 -255
rect 388 -451 444 -441
rect 388 -765 444 -755
rect 388 -951 444 -941
rect 142 -1265 198 -1255
rect 142 -1451 198 -1441
rect 302 -1265 354 -1255
rect 302 -1451 354 -1441
rect 311 -1553 345 -1451
rect -5 -1584 345 -1553
<< via2 >>
rect -104 59 -102 235
rect -102 59 -50 235
rect -50 59 -48 235
rect 142 59 144 235
rect 144 59 196 235
rect 196 59 198 235
rect 142 -441 144 -265
rect 144 -441 196 -265
rect 196 -441 198 -265
rect 142 -941 144 -765
rect 144 -941 196 -765
rect 196 -941 198 -765
rect -104 -1441 -102 -1265
rect -102 -1441 -50 -1265
rect -50 -1441 -48 -1265
rect 388 -441 390 -265
rect 390 -441 442 -265
rect 442 -441 444 -265
rect 388 -941 390 -765
rect 390 -941 442 -765
rect 442 -941 444 -765
rect 142 -1441 144 -1265
rect 144 -1441 196 -1265
rect 196 -1441 198 -1265
<< metal3 >>
rect -114 380 454 440
rect -114 235 -38 380
rect -114 59 -104 235
rect -48 59 -38 235
rect -114 -1265 -38 59
rect -114 -1441 -104 -1265
rect -48 -1441 -38 -1265
rect -114 -1586 -38 -1441
rect 132 235 208 240
rect 132 59 142 235
rect 198 59 208 235
rect 132 -265 208 59
rect 132 -441 142 -265
rect 198 -441 208 -265
rect 132 -765 208 -441
rect 132 -941 142 -765
rect 198 -941 208 -765
rect 132 -1265 208 -941
rect 132 -1441 142 -1265
rect 198 -1441 208 -1265
rect 132 -1446 208 -1441
rect 378 -265 454 380
rect 378 -441 388 -265
rect 444 -441 454 -265
rect 378 -765 454 -441
rect 378 -941 388 -765
rect 444 -941 454 -765
rect 378 -1586 454 -941
rect -114 -1646 454 -1586
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729246161
transform 1 0 -32 0 1 147
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729246161
transform 1 0 372 0 1 -853
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729246161
transform 1 0 372 0 1 147
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729246161
transform 1 0 -32 0 1 -353
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729246161
transform 1 0 372 0 1 -353
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729246161
transform 1 0 -32 0 1 -853
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729246161
transform 1 0 -32 0 1 -1353
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729246161
transform 1 0 372 0 1 -1353
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729246161
transform 1 0 170 0 1 -1353
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729246161
transform 1 0 170 0 1 147
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_2
timestamp 1729246161
transform 1 0 170 0 1 -353
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_3
timestamp 1729246161
transform 1 0 170 0 1 -853
box -223 -200 223 200
<< labels >>
flabel viali 91 482 91 482 0 FreeSans 480 0 0 0 vdd
port 0 nsew
flabel metal2 327 361 327 361 0 FreeSans 480 0 0 0 d6
port 1 nsew
flabel via2 -76 -1354 -76 -1354 0 FreeSans 480 0 0 0 out
port 3 nsew
flabel via1 249 -1189 249 -1189 0 FreeSans 480 0 0 0 vin
port 4 nsew
flabel metal1 91 -68 91 -68 0 FreeSans 480 0 0 0 vip
port 5 nsew
flabel metal3 169 -609 169 -609 0 FreeSans 480 0 0 0 d5
port 6 nsew
<< end >>
