magic
tech sky130A
magscale 1 2
timestamp 1729183514
<< pwell >>
rect -840 -737 840 737
<< nmos >>
rect -644 -527 644 527
<< ndiff >>
rect -702 515 -644 527
rect -702 -515 -690 515
rect -656 -515 -644 515
rect -702 -527 -644 -515
rect 644 515 702 527
rect 644 -515 656 515
rect 690 -515 702 515
rect 644 -527 702 -515
<< ndiffc >>
rect -690 -515 -656 515
rect 656 -515 690 515
<< psubdiff >>
rect -804 667 -708 701
rect 708 667 804 701
rect -804 605 -770 667
rect 770 605 804 667
rect -804 -667 -770 -605
rect 770 -667 804 -605
rect -804 -701 -708 -667
rect 708 -701 804 -667
<< psubdiffcont >>
rect -708 667 708 701
rect -804 -605 -770 605
rect 770 -605 804 605
rect -708 -701 708 -667
<< poly >>
rect -644 599 644 615
rect -644 565 -628 599
rect 628 565 644 599
rect -644 527 644 565
rect -644 -565 644 -527
rect -644 -599 -628 -565
rect 628 -599 644 -565
rect -644 -615 644 -599
<< polycont >>
rect -628 565 628 599
rect -628 -599 628 -565
<< locali >>
rect -804 667 -708 701
rect 708 667 804 701
rect -804 605 -770 667
rect 770 605 804 667
rect -644 565 -628 599
rect 628 565 644 599
rect -690 515 -656 531
rect -690 -531 -656 -515
rect 656 515 690 531
rect 656 -531 690 -515
rect -644 -599 -628 -565
rect 628 -599 644 -565
rect -804 -667 -770 -605
rect 770 -667 804 -605
rect -804 -701 -708 -667
rect 708 -701 804 -667
<< viali >>
rect -628 565 628 599
rect -690 -515 -656 515
rect 656 -515 690 515
rect -628 -599 628 -565
<< metal1 >>
rect -640 599 640 605
rect -640 565 -628 599
rect 628 565 640 599
rect -640 559 640 565
rect -696 515 -650 527
rect -696 -515 -690 515
rect -656 -515 -650 515
rect -696 -527 -650 -515
rect 650 515 696 527
rect 650 -515 656 515
rect 690 -515 696 515
rect 650 -527 696 -515
rect -640 -565 640 -559
rect -640 -599 -628 -565
rect 628 -599 640 -565
rect -640 -605 640 -599
<< properties >>
string FIXED_BBOX -787 -684 787 684
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.27 l 6.44 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
